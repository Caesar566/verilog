module JK_trigger (
    
);

endmodule //JK_trigger